--------------------------------------------------------------------------------
-- Title       : <Title Block>
-- Project     : Default Project Name
--------------------------------------------------------------------------------
-- File        : Filtro_Digital_tb.vhd
-- Author      : User Name <user.email@user.company.com>
-- Company     : User Company Name
-- Created     : Mon May 17 14:30:31 2021
-- Last update : Mon May 17 14:30:31 2021
-- Platform    : Default Part Number
-- Standard    : <VHDL-2008 | VHDL-2002 | VHDL-1993 | VHDL-1987>
--------------------------------------------------------------------------------
-- Copyright (c) 2021 User Company Name
-------------------------------------------------------------------------------
-- Description: 
--------------------------------------------------------------------------------
-- Revisions:  Revisions and documentation are controlled by
-- the revision control system (RCS).  The RCS should be consulted
-- on revision history.
-------------------------------------------------------------------------------

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use std.textio.all;
use ieee.std_logic_textio.all;

-----------------------------------------------------------

entity Filtro_Digital_tb is

end entity Filtro_Digital_tb;

-----------------------------------------------------------

architecture testbench of Filtro_Digital_tb is

	-- Testbench DUT generics


	-- Testbench DUT ports
	signal clk     : std_logic;
	signal rst     : std_logic;
	signal CHA     : std_logic;
	signal CHB     : std_logic;
	signal CHA_out : std_logic;
	signal CHB_out : std_logic;

	-- Other constants
	constant C_CLK_PERIOD : real := 10.0e-9; -- NS

begin
	-----------------------------------------------------------
	-- Clocks and Reset
	-----------------------------------------------------------
	CLK_GEN : process
	begin
		clk <= '1';
		wait for C_CLK_PERIOD / 2.0 * (1 SEC);
		clk <= '0';
		wait for C_CLK_PERIOD / 2.0 * (1 SEC);
	end process CLK_GEN;

   -- process
	--begin
		--CHA <= '1';
		--wait for 1 ms;
		--CHB <= '1';
		--wait for 3 ms;
		--CHA <= '0';
		--wait for 1 ms;
		--CHB <= '0';
		--wait for 3 ms;
	--end process;


	RESET_GEN : process
	begin
		rst <= '1';
		CHA <= '0';
		CHB <= '0';
		wait for 3 us;
		rst <= '0';
		CHA <= '1';
		wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';

        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 ns;
        CHB <= '0';
        wait for 3 ns;
        CHA <= '1';
        wait for 1 ns;
        CHB <= '1';
        wait for 3 ns;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
        wait for 3 us;
        CHA <= '0';
        wait for 1 us;
        CHB <= '0';
        wait for 3 us;
        CHA <= '1';
        wait for 1 us;
		CHB <= '1';
		


        
		wait;
	end process RESET_GEN;

	-----------------------------------------------------------
	-- Testbench Stimulus
	-----------------------------------------------------------

	-----------------------------------------------------------
	-- Entity Under Test
	-----------------------------------------------------------
	DUT : entity work.Filtro_Digital
		port map (
			clk     => clk,
			rst     => rst,
			CHA     => CHA,
			CHB     => CHB,
			CHA_out => CHA_out,
			CHB_out => CHB_out
		);

end architecture testbench;